-- uart_tx_fsm.vhd: UART controller - finite state machine controlling TX side
-- Author(s): Name Surname (xlogin00)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;



entity UART_TX_FSM is
    port(
       CLK : in std_logic;
       RST : in std_logic
    );
end entity;



architecture behavioral of UART_TX_FSM is
begin

end architecture;
